module program_counter(input clk, rst, take_branch, take_jump, take_jr, input [31:0] branch_offset, input [25:0] jump_offset, input [31:0] jr_addr, output reg [31:0] pc);
    
    
endmodule